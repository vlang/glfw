module main

fn main() {

}
